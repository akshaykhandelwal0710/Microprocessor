module control_signal_decoder #(parameter sz = 20, parameter SZ = 24)(
  input [sz-1:0] val_in,
  output [SZ-1:0] val_out
);
  
endmodule